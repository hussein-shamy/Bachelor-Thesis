//////////////////////////////////////////////////////////////////////////////////
//	
//								Tanta University
//						   	 Faculty of Engineering
//		Electronics and Electrical Communications Engineering Department
//
//////////////////////////////////////////////////////////////////////////////////
//
// Project Name: 	Meeting 5G Latency Requirements in Cell Outage Compensation (COC) 
//               	in Self Organizing Networks (SONs) using Hardware Acceleration.
//
// Create Date:    03/Feb/2023 
// Module Name:    PRNG 
// Design Name:    Q_Learining_SON
// Engineers:	   Mohamed Hellal
//
//////////////////////////////////////////////////////////////////////////////////
//discription:
// The PRNG module is a simple pseudorandom number generator (PRNG) based on a linear feedback shift register (LFSR) architecture.
// It generates a 16-bit PRNG output, PRNG_out, and provides the Action output as the two most significant bits of PRNG_out.
// The module has inputs CLK and RST for clocking and resetting the PRNG.
// The module includes a register, PRNG_out, to store the PRNG output.
// The feedback signal is generated by XORing the last two bits (bit 15 and bit 13) and two additional bits (bits 12 and 10) of PRNG_out.
// The Action output is assigned the two most significant bits (bits 13 and 12) of PRNG_out.
// The module uses a synchronous always block with posedge CLK and negedge RST to generate the PRNG output.
// When not in reset, the module shifts the PRNG_out left by one bit and appends the feedback bit to the LSB position.
// The initial value of PRNG_out is set to the Seed value during reset.
//////////////////////////////////////////////////////////////////////////////////


module PRNG #(parameter Seed = 16'b1000001000101000) (
  input 	wire CLK, RST,       	// Clock and Reset signals
  output 	reg	 [3:0] Action   	// Output signal representing the two most significant bits of PRNG_out
);

  reg [15:0] PRNG_out;       // Register to store the PRNG output
  wire feedback;             // Feedback signal for XORing the last two bits of PRNG_out
	
//feedback is XORing the 15,13,12,10
assign feedback = PRNG_out[15] ^ PRNG_out[13] ^ PRNG_out[12] ^ PRNG_out[10];

//assign action the two MSBs from PRNG_out
// assign	Action = PRNG_out[15:12];

//  main PRNG code

always @(posedge CLK, negedge RST)
begin
 if (!RST)
 begin
	PRNG_out <= Seed;                                // Reset PRNG_out to the predefined Seed value
 end
 else
 begin
	PRNG_out[15:0] <= {PRNG_out[14:0], feedback};    // Shift PRNG_out left by one bit and append the feedback bit
 end
end

//RandomNum - Action mapping
always@(*)
begin
	case (PRNG_out[15:12])
	4'b0000:	Action = 4'b0000;
	4'b0001:	Action = 4'b0000;
	4'b0010:	Action = 4'b0001;
	4'b0011:	Action = 4'b0001;
	4'b0100:	Action = 4'b0010;
	4'b0101:	Action = 4'b0010;
	4'b0110:	Action = 4'b0011;
	4'b0111:	Action = 4'b0011;
	4'b1000:	Action = 4'b0100;
	4'b1001:	Action = 4'b0100;
	4'b1010:	Action = 4'b0101;
	4'b1011:	Action = 4'b0101;
	4'b1100:	Action = 4'b0110;
	4'b1101:	Action = 4'b0110;
	4'b1110:	Action = 4'b0111;
	4'b1111:	Action = 4'b1000;
endcase
end

endmodule