`timescale 1us/1ns
module PQL_TOP_tb ();

reg					CLK,RST;
reg		[95:0]		RS0,RS1,RS2,RS3,RS4,RS5;
reg		[23:0]		alpha, Gamma;

wire	[23:0]		Q0_0	,Q0_1	,Q0_2	,Q0_3,    	// from Sn with parameter (state_num = 0)
					Q1_0	,Q1_1	,Q1_2	,Q1_3,    	// from Sn with parameter (state_num = 1)
					Q2_0	,Q2_1	,Q2_2	,Q2_3,    	// from Sn with parameter (state_num = 2)
					Q3_0	,Q3_1	,Q3_2	,Q3_3,    	// from Sn with parameter (state_num = 3)
					Q4_0	,Q4_1	,Q4_2	,Q4_3,    	// from Sn with parameter (state_num = 4)
                    Q5_0	,Q5_1	,Q5_2	,Q5_3;					// from Sn with parameter (state_num = 5)
					
PQL_Top DUT (
.CLK    (CLK),
.RST    (RST),
.RS0    (RS0),
.RS1    (RS1),
.RS2    (RS2),
.RS3    (RS3),
.RS4    (RS4),
.RS5    (RS5),
.alpha	(alpha),
.Gamma	(Gamma),
.Q0_0(Q0_0)	,.Q0_1(Q0_1)	,.Q0_2(Q0_2)	,.Q0_3(Q0_3),
.Q1_0(Q1_0)	,.Q1_1(Q1_1)	,.Q1_2(Q1_2)	,.Q1_3(Q1_3),
.Q2_0(Q2_0)	,.Q2_1(Q2_1)	,.Q2_2(Q2_2)	,.Q2_3(Q2_3),
.Q3_0(Q3_0)	,.Q3_1(Q3_1)	,.Q3_2(Q3_2)	,.Q3_3(Q3_3),
.Q4_0(Q4_0)	,.Q4_1(Q4_1)	,.Q4_2(Q4_2)	,.Q4_3(Q4_3),
.Q5_0(Q5_0)	,.Q5_1(Q5_1)	,.Q5_2(Q5_2)	,.Q5_3(Q5_3)
);

initial begin
	$dumpfile("PQL_TOP_tb_14.vcd");
	$dumpvars;
	
	CLK     = 0;
	RST     = 1;
	RS0     = 96'b000000000000000000000000_111111010000000000000000_000000000000000000000000_111111010000000000000000;
	RS1     = 96'b000000000000000000000000_000000000000000000000000_000000000000000000000000_111111010000000000000000;
	RS2     = 96'b111111010000000000000000_000000000000000000000000_000110010000000000000000_111111010000000000000000;
	RS3     = 96'b000000000000000000000000_111111010000000000000000_111111010000000000000000_000000000000000000000000;
	RS4     = 96'b000110010000000000000000_000000000000000000000000_111111010000000000000000_000000000000000000000000;
	RS5     = 96'b111111010000000000000000_000000000000000000000000_111111010000000000000000_000000000000000000000000;
	alpha   = 24'b0000000000011001100110011;
	Gamma	= 24'b0000000000011001100110011;
	
	#1;
	RST = 0;
	#1;
	RST = 1;
	
	#640000;
	$stop;
end

always #5 CLK=~CLK;

endmodule